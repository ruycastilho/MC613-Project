LIBRARY ieee ; 
USE ieee.std_logic_1164.all;
LIBRARY work; 
USE work.data_types.all;

ENTITY serial IS 
	PORT (
			image:		IN image_array);

END serial;

ARCHITECTURE Behavior OF serial IS
	BEGIN

				
END Behavior ;